* Prova SEL0622 - Questao 10 - Simulacao sobre layout do circuito contador
*                              com opcao de extracao R+C+CC
*
* entradas: 
*       - CLK   : Pulso de clock de entrada
*       - RESET : Sincrono e volta a contagem para zero
*
* saidas:
*       - COUNT1(4 downto 0) : valor binario da contagem
*       - CLKDIV : pulso dividido por 29
*
* @author: Rodrigo Ferrari
* @date: 11/01/18
.option list
.defmod NMOS4 MODN
.defmod PMOS4 MODP

* Usar modelo tipico de simulacao 'tm';
* outros modelos: 'wp' e 'ws'
.lib "/local/tools/dkit/ams_3.70_mgc/eldo/c35/wc53.lib" tm

* Importar netlists e verificar ordem da definicao do subcircuito
.include "../../cu.lib/default.group/layout.views/contador/contador.cal/contador.pex.netlist"
Xcont RESET CLK COUNT1[0] COUNT1[2] COUNT1[4] COUNT1[3] COUNT1[1] VDD VSS CONTADOR

.param vd=3v
.param F1='0.5G'
.param T1='1/F1'
.param TDEL='0.1*T1'

* tempo de simul
.param ST='120*T1'
.param STEP='0.5*T1'

* circuito
.connect VSS 0
.connect RESET VSS
.connect CLKDIV COUNT1[4]
VDD_S VDD VSS vd
Vclk CLK VSS PULSE(0 3 0 TDEL TDEL 'T1/2 - TDEL' T1)

.op
.tran 1 ST 0 STEP sweep F1 0.45G 0.60G  0.01G
*.tran 1 ST 0 STEP
.plot tran V(CLK) V(COUNT1[0]) V(COUNT1[1]) V(COUNT1[2]) V(COUNT1[3]) V(COUNT1[4]) V(CLKDIV)

* medidas
.meas tran ti trig V(CLK)    val='vd/2' fall=50 targ v(CLK)    val='vd/2' fall=51
.meas tran to trig V(CLKDIV) val='vd/2' fall=2  targ V(CLKDIV) val='vd/2' fall=3
.meas tran fi param='1/ti'
.meas tran fo param='1/to'
.meas tran div param='fi/fo'
.meas tran iavg avg Is(vdd_s)
.meas tran power param='-iavg*vd'
.meas tran cons param='((power/(1m))/(F1/(1G)))'
.end
